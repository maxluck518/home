always @(posedge clk) begin
    if (!reset) begin
    end
    else begin
    end
end
