module inst3(/*vlog_aide:auto_port*/);

input           inst3_in0;
input [5:0]     inst3_in1;
output [7:0]    inst3_out0;

endmodule
