module auto_port(/*vlog_aide:auto_port*/);

input           test1;
input           test21, test22, test23;
input [3:0]     test3;
input [`DATA_WIDTH-1:0] test4;
output          test5, test51;
output  [15:0]  test6;
inout           test7;

endmodule
