interface  ();
// Input ports of DUT
logic [ 3:0] IMP_SEL_FS;
logic  PD18_VDDR_G;
logic [7:0] RESERVE_IN;
logic  VG_IN_PHASE;
logic  VBUS_ON;
// Output ports of DUT
logic  VG_OUT_PHASE;
logic  PD18_VDDR_G_OUT;
logic [7:0] RESERVE_OUT;
// Inout ports of DUT
endinterface
